// Code your design here
module not_struc(a,y);
  input a;
  output y;
  not g1(y,a);
endmodule
